0: mdr = {`LOAD, 5'd13};
1: mdr = {`STORE, 5'd16};
2: mdr = {`LOAD, 5'd14};
3: mdr = {`STORE, 5'd17};
4: mdr = {`STORE, 5'd31};
5: mdr = {`LOAD, 5'd16};
6: mdr = {`ADD, 5'd17};
7: mdr = {`STORE, 5'd18};
8: mdr = {`LOAD, 5'd17};
9: mdr = {`STORE, 5'd16};
10: mdr = {`LOAD, 5'd18};
11: mdr = {`STORE, 5'd17};
12: mdr = {`BNE, 5'd15};
13: mdr = {`LOAD, 5'd0};
14: mdr = {`LOAD, 5'd1};
15: mdr = {`LOAD, 5'd5};
