0: mdr = {`LOAD, 5'd13};
1: mdr = {`STORE, 5'd16};
2: mdr = {`STORE, 5'd17};
3: mdr = {`STORE, 5'd31};
4: mdr = {`LOAD, 5'd16};
5: mdr = {`ADD, 5'd17};
6: mdr = {`STORE, 5'd18};
7: mdr = {`STORE, 5'd31};
8: mdr = {`LOAD, 5'd17};
9: mdr = {`STORE, 5'd16};
10: mdr = {`LOAD, 5'd18};
11: mdr = {`STORE, 5'd17};
12: mdr = {`BNE, 5'd14};
13: mdr = {`LOAD, 5'd1};
14: mdr = {`LOAD, 5'd4};
